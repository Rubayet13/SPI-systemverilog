package env_pkg;

  import agent_pkg::*;

  `include "spi_sco.sv"
  `include "spi_env.sv"

endpackage