package agent_pkg;

    `include "spi_trans.sv"
    `include "spi_driver.sv"
    `include "spi_monitor.sv"
    `include "spi_generator.sv"
    
endpackage